module test(a, b);
	input [5:0] a;
	output [5:0] b;
	assign b[0] = 1;
	assign b[1] = 0;
	assign b[2] = 0;
	assign b[3] = 0;
	assign b[4] = 0;
	assign b[5] = 0;
endmodule